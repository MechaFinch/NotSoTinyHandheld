--
-- Mechafinch
-- NST Handheld Project
-- 
-- nst_instruction_cache
-- Instruction cache.
-- 2-way set associative, LRU, read only
-- 256 sets with 8 byte blocks
-- Uses 9 BRAM blocks
--

library ieee;
use ieee.std_logic_1164.all;
use work.nst_types.all;

library efxphysicallib;
use efxphysicallib.efxcomponents.all;

entity nst_insturction_cache is
	port (
		-- cpu side
		address:	in nst_dword_t;				-- address the cpu is reading
		data:		out icache_block_data_t;	-- data block for the cpu
		data_ready:	out std_logic;
		
		-- memory side
		mem_address:	out nst_dword_t;		-- address the cache is reading
		mem_data:		in icache_block_data_t;	-- data block for the cache
		mem_ready:		in std_logic;
		
		-- clocking
		exec_clk:	in std_logic;
	);
end nst_instruction_cache;

architecture a1 of nst_instruction_cache is
	-- a block; data with tag and dirty bit
	type icache_block_t is record
		data: 	icache_block_data_t; -- array of 8 bytes
		tag:	std_logic_vector(20 downto 0);
		clean:	std_logic; -- 0 = dirty, for ease of initialization
	end record;
	
	-- a set; 2 blocks with LRU and valid bits
	-- There is only one valid bit per set in order to save a BRAM (in doing so not wasting 90% of one)
	-- When data is read into an invalid set, it is written to both blocks (they recieve the same tag)
	-- to prevent false hits. When both blocks in a set match an address, b0 will be used. 
	type icache_set_t is record
		b0:		icache_block_t;
		b1:		icache_block_t;
		lru:	std_logic;	-- 0 = b0 LRU, 1 = b1 LRU
		valid:	std_logic;	-- 0 = invalid, 1 = valid
	end record;
	
	type bram_data_t is array (8 downto 0) of std_logic_vector(19 downto 0);
	
	signal current_input:	icache_set_t;
	signal current_output:	icache_set_t;
	
	signal bram_write_enable:	std_logic;
	signal bram_address:		std_logic_vector(11 downto 0);
	
	signal bram_inputs:		bram_data_t;
	signal bram_outputs:	bram_data_t;
begin

	-- BRAM address is the set index subset of the address
	bram_addr_proc: process (all) begin
		-- only the upper 8 bits of address are used
		-- primitives doc says to leave lines not used by the mode unconnected
		bram_address(11 downto 4)	<= address(10 downto 3);
		bram_address(3 downto 0)	<= open;
	end process;
	
	-- handles renaming input/output as a cache set record and as bram signals
	bram_mapping_proc: process (all) begin
		-- BRAM input mapping
		-- block 0: bits 19:0 of b0; bits 19:0 of b0's data
		bram_inputs(0)(7 downto 0)		<= current_input.b0.data(0);
		bram_inputs(0)(15 downto 8)		<= current_input.b0.data(1);
		bram_inputs(0)(19 downto 16)	<= current_input.b0.data(2)(3 downto 0);
		
		-- block 1: bits 39:20 of b0; bits 39:20 of b0's data
		bram_inputs(1)(3 downto 0)		<= current_input.b0.data(2)(7 downto 4);
		bram_inputs(1)(11 downto 4)		<= current_input.b0.data(3);
		bram_inputs(1)(19 downto 12)	<= current_input.b0.data(4);
		
		-- block 2: bits 59:40 of b0; bits 59:40 of b0's data
		bram_inputs(2)(7 downto 0)		<= current_input.b0.data(5);
		bram_inputs(2)(15 downto 8)		<= current_input.b0.data(6);
		bram_inputs(2)(19 downto 16)	<= current_input.b0.data(7)(3 downto 0);
		
		-- block 3: bits 79:60 of b0; bits 63:60 of b0's data, 15:0 of b0's tag
		bram_inputs(3)(3 downto 0)	<= current_input.b0.data(7)(7 downto 4);
		bram_inputs(3)(19 downto 4)	<= current_input.b0.tag(15 downto 0);
		
		-- block 4: bits 85:80 of b0, 7:0 of b1; bits 20:16 of b0's tag, b0's clean bit, bits 7:0 of b1's data
		bram_inputs(4)(4 downto 0)		<= current_input.b0.tag(20 downto 16);
		bram_inputs(4)(5)				<= current_input.b0.clean;
		bram_inputs(4)(11 downto 6)		<= "000000"; -- 6 unused bits, aligns very conveniently
		bram_inputs(4)(19 downto 12)	<= current_input.b1.data(0);
		
		-- block 5: bits 27:8 of b1; bits 27:8 of b1's data
		bram_inputs(5)(7 downto 0)		<= current_input.b1.data(1);
		bram_inputs(5)(15 downto 8)		<= current_input.b1.data(2);
		bram_inputs(5)(19 downto 16)	<= current_input.b1.data(3)(3 downto 0);
		
		-- block 6: bits 47:28 of b1; bits 47:28 of b1's data
		bram_inputs(6)(3 downto 0)		<= current_input.b1.data(3)(7 downto 4);
		bram_inputs(6)(11 downto 4)		<= current_input.b1.data(4);
		bram_inputs(6)(19 downto 12)	<= current_input.b1.data(5);
		
		-- block 7: bits 67:48 of b1; bits 63:48 of b1's data, 3:0 of b1's tag
		bram_inputs(7)(7 downto 0)		<= current_input.b1.data(6);
		bram_inputs(7)(15 downto 8)		<= current_input.b1.data(7);
		bram_inputs(7)(19 downto 16)	<= current_input.b1.tag(3 downto 0);
		
		-- block 8: bits 85:68 of b1, set status bits; bits 20:4 of b1's tag, b1's clean bit, set LRU bit, set valid bit
		bram_inputs(8)(16 downto 0)	<= current_input.b1.tag(20 downto 4);
		bram_inputs(8)(17)			<= current_input.b1.clean;
		bram_inputs(8)(18)			<= current_input.lru;
		bram_inputs(8)(19)			<= current_input.valid;
		
		-- BRAM output mapping (see above)
		current_output.b0.data(0)				<= bram_outputs(0)(7 downto 0);
		current_output.b0.data(1)				<= bram_outputs(0)(15 downto 8);
		current_output.b0.data(2)(7 downto 4)	<= bram_outputs(1)(3 downto 0);
		current_output.b0.data(2)(3 downto 0)	<= bram_outputs(0)(19 downto 16);
		current_output.b0.data(3)				<= bram_outputs(1)(11 downto 4);
		current_output.b0.data(4)				<= bram_outputs(1)(19 downto 12);
		current_output.b0.data(5)				<= bram_outputs(2)(7 downto 0);
		current_output.b0.data(6)				<= bram_outputs(2)(15 downto 8);
		current_output.b0.data(7)(7 downto 4)	<= bram_outputs(3)(3 downto 0);
		current_output.b0.data(7)(3 downto 0)	<= bram_outputs(2)(19 downto 16);
		
		current_output.b0.tag(20 downto 16)	<= bram_outputs(4)(4 downto 0);
		current_output.b0.tag(15 downto 0)	<= bram_outputs(3)(19 downto 4);
		current_output.b0.clean				<= bram_outputs(4)(5);
		
		current_output.b1.data(0)				<= bram_outputs(4)(19 downto 12);
		current_output.b1.data(1)				<= bram_outputs(5)(7 downto 0);
		current_output.b1.data(2)				<= bram_outputs(5)(15 downto 8);
		current_output.b1.data(3)(7 downto 4)	<= bram_outputs(6)(3 downto 0);
		current_output.b1.data(3)(3 downto 0)	<= bram_outputs(5)(19 downto 16);
		current_output.b1.data(4)				<= bram_outputs(6)(11 downto 4);
		current_output.b1.data(5)				<= bram_outputs(6)(19 downto 12);
		current_output.b1.data(6)				<= bram_outputs(7)(7 downto 0);
		current_output.b1.data(7)				<= bram_outputs(7)(15 downto 8);
		
		current_output.b1.tag(20 downto 4)	<= bram_outputs(8)(16 downto 0);
		current_output.b1.tag(3 downto 0)	<= bram_outputs(7)(19 downto 16);
		current_output.b1.clean				<= bram_outputs(8)(17);
		
		current_output.lru		<= bram_outputs(8)(18);
		current_output.valid	<= bram_outputs(8)(19);
	end process;

	-- BRAM instances
	-- Each BRAM is addressed by the set number
	
	-- block 0: bits 19:0 of the set; bits 19:0 of b0; bits 19:0 of b0's data
	bram_0: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(0),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(0)
		);
	
	-- block 1: bits 39:20 of the set; bits 39:20 of b0; bits 39:20 of b0's data
	bram_1: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(1),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(1)
		);
		
	-- block 2: bits 59:40 of the set; bits 59:40 of b0; bits 59:40 of b0's data
	bram_2: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(2),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(2)
		);
		
	-- block 3: bits 79:60 of the set; bits 79:60 of b0; bits 63:60 of b0's data, 15:0 of b0's tag
	bram_3: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(3),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(3)
		);
		
	-- block 4: bits 99:80 of the set; bits 85:80 of b0, 13:0 of b1; bits 20:16 of b0's tag, b0's clean bit, bits 13:0 of b1's data
	bram_4: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(4),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(4)
		);
		
	-- block 5: bits 119:100 of the set; bits 33:14 of b1; bits 33:14 of b1's data
	bram_5: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(5),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(5)
		);
		
	-- block 6: bits 139:120 of the set; bits 53:34 of b1; bits 53:34 of b1's data
	bram_6: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(6),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(6)
		);
		
	-- block 7: bits 159:140 of the set; bits 73:54 of b1; bits 63:54 of b1's data, 9:0 of b1's tag
	bram_7: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(7),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(7)
		);
		
	-- block 8: bits 173:160 of the set; bits 85:74 of b1, set status bits; bits 20:10 of b1's tag, b1's clean bit, set LRU bit, set valid bit
	bram_8: EFX_RAM_5K
		generic map (
			READ_WIDTH	=> 20,
			WRITE_WIDTH	=> 20,
			OUTPUT_REG	=> '0',
			WRITE_MODE	=> "READ_UNKNOWN", 
			
			WCLK_POLARITY	=> '1',	-- rising edge
			WCLKE_POLARITY	=> '1',
			WE_POLARITY		=> '1',
			
			RCLK_POLARITY	=> '0',	-- falling edge
			RE_POLARITY		=> '1',
		
			INIT_0	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_1	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_2	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_3	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_4	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_5	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_6	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_7	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_8	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_9	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_A	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_B	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_C	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_D	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_E	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_F	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_10	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_11	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_12	=> 256x"0000000000000000000000000000000000000000000000000000000000000000",
			INIT_13	=> 256x"0000000000000000000000000000000000000000000000000000000000000000"
		)
		port map (
			WCLK	=> exec_clk,
			WE		=> bram_write_enable,
			WCLKE	=> '1',
			RCLK	=> exec_clk,
			RE		=> '1',
			WADDR	=> bram_address,
			WDATA	=> bram_outputs(8),
			RADDR	=> bram_address,
			RDATA	=> bram_inputs(8)
		);
		
	
	
end a1;