--
-- Mechafinch
-- NST Handheld Project
--
-- nst_control
-- Control logic for the CPU. A lot of this is a big ole lookup table from the (converted) opcode
-- to most of the control signals.
--
