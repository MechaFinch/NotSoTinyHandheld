--
-- Mechafinch
-- NST Handheld Project
--
-- nst_spi_interface
-- SPI bus interface. This module will operate the SPI bus, including interrupts, memory-mapped
-- IO/config, and so on.
--